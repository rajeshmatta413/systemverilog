// -------------------------------------------------------
// -- hi
// -------------------------------------------------------
